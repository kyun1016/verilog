`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:15:08 10/18/2019 
// Design Name: 
// Module Name:    my_application 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module my_application(
    input clk,
    input A,
    input B,
    output [3:0] num,
    output state
    );


//�������¸� �����ϴ� ����ȸ�� ���

//������¸� �����ϴ� ����ȸ�� ���

//��°��� �����ϴ� ����ȸ�� ���

endmodule
